--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:36:27 02/10/2016
-- Design Name:   
-- Module Name:   /home/craig/Documents/Projects/Repos/OT_1588_Master/OT_1588_Master/TB_nmea_lcd_display_ctrl.vhd
-- Project Name:  vault_numato
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: nmea_lcd_display_ctrl
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY TB_nmea_lcd_display_ctrl IS
END TB_nmea_lcd_display_ctrl;
 
ARCHITECTURE behavior OF TB_nmea_lcd_display_ctrl IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT nmea_lcd_display_ctrl
    PORT(
         CLK_IN : IN  std_logic;
         RST_IN : IN  std_logic;
         ADDR_OUT : OUT  std_logic_vector(7 downto 0);
         DATA_IN : IN  std_logic_vector(7 downto 0);
         LINE1_OUT : OUT  std_logic_vector(127 downto 0);
         LINE2_OUT : OUT  std_logic_vector(127 downto 0)
        );
    END COMPONENT;

    COMPONENT nmea_parser
    PORT(
         CLK_IN         : IN  std_logic;
         RST_IN         : IN  std_logic;
         NMEA_EN_IN     : IN  std_logic;
         NMEA_DATA_IN   : IN  std_logic_vector(7 downto 0);
         ADDR_IN        : IN  std_logic_vector(7 downto 0);
         DATA_OUT       : OUT  std_logic_vector(7 downto 0));
    END COMPONENT;

   --Inputs
   signal CLK_IN : std_logic := '0';
   signal RST_IN : std_logic := '0';
   signal DATA_IN : std_logic_vector(7 downto 0) := (others => '0');

   signal NMEA_EN_IN    : std_logic := '0';
   signal NMEA_DATA_IN  : std_logic_vector(7 downto 0) := (others => '0');

 	--Outputs
   signal ADDR_OUT : std_logic_vector(7 downto 0);
   signal LINE1_OUT : std_logic_vector(127 downto 0);
   signal LINE2_OUT : std_logic_vector(127 downto 0);

   -- Clock period definitions
   constant CLK_IN_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: nmea_lcd_display_ctrl PORT MAP (
          CLK_IN => CLK_IN,
          RST_IN => RST_IN,
          ADDR_OUT => ADDR_OUT,
          DATA_IN => DATA_IN,
          LINE1_OUT => LINE1_OUT,
          LINE2_OUT => LINE2_OUT
        );

   uut2: nmea_parser PORT MAP (
          CLK_IN        => CLK_IN,
          RST_IN        => RST_IN,
          NMEA_EN_IN    => NMEA_EN_IN,
          NMEA_DATA_IN  => NMEA_DATA_IN,
          ADDR_IN       => ADDR_OUT,
          DATA_OUT      => DATA_IN
        );

   -- Clock process definitions
   CLK_IN_process :process
   begin
		CLK_IN <= '0';
		wait for CLK_IN_period/2;
		CLK_IN <= '1';
		wait for CLK_IN_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for CLK_IN_period * 1000;  

      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"56";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4b";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"52";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"43";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"56";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4b";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"52";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"43";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"56";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4b";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"46";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"52";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"43";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"56";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4b";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"56";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"56";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"56";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"52";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"43";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"56";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4b";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"44";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"52";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"43";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"56";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4b";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"43";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"52";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"43";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"53";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"35";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"38";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"45";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"32";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"31";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"36";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"37";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"24";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"50";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"56";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"47";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"33";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"34";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"39";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"54";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4d";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2e";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"4b";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2c";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"2a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"30";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"41";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;
      NMEA_EN_IN <= '1';
      NMEA_DATA_IN <= X"0a";
      wait for CLK_IN_period;
      NMEA_EN_IN <= '0';
      wait for CLK_IN_period * 20;

      wait;
   end process;

END;
