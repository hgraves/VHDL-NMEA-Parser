--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   15:05:13 02/09/2016
-- Design Name:   
-- Module Name:   /home/craig/Documents/Projects/Repos/OT_1588_Master/OT_1588_Master/TB_nmea_parser.vhd
-- Project Name:  vault_numato
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: nmea_parser
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY TB_nmea_parser IS
END TB_nmea_parser;
 
ARCHITECTURE behavior OF TB_nmea_parser IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT nmea_parser
    PORT(
         CLK_IN         			: IN  std_logic;
         RST_IN         			: IN  std_logic;
         NMEA_EN_IN     			: IN  std_logic;
         NMEA_DATA_IN   			: IN  std_logic_vector(7 downto 0);
         NMEA_EN_OUT    			: OUT STD_LOGIC;
         NMEA_DATA_OUT  			: OUT STD_LOGIC_VECTOR(7 downto 0);
         NMEA_EN_ACK_IN 			: IN STD_LOGIC;
			NEW_TIMESTAMP_EN_OUT    : OUT STD_LOGIC;
         TIMESTAMP_DATA_OUT      : OUT STD_LOGIC_VECTOR(31 downto 0);
         ADDR_IN        			: IN  std_logic_vector(7 downto 0);
         DATA_OUT       			: OUT  std_logic_vector(7 downto 0));
    END COMPONENT;
    
    COMPONENT uart
    generic (
        baud                : positive;
        clock_frequency     : positive
    );
    port (  
        clock               :   in  std_logic;
        reset               :   in  std_logic;    
        data_stream_in      :   in  std_logic_vector(7 downto 0);
        data_stream_in_stb  :   in  std_logic;
        data_stream_in_ack  :   out std_logic;
        data_stream_out     :   out std_logic_vector(7 downto 0);
        data_stream_out_stb :   out std_logic;
        tx                  :   out std_logic;
        rx                  :   in  std_logic
    );
    END COMPONENT;

   --Inputs
   signal CLK_IN        			: std_logic := '0';
   signal RST_IN        			: std_logic := '0';
   signal NMEA_EN_IN    			: std_logic := '0';
   signal NMEA_DATA_IN  			: std_logic_vector(7 downto 0) := (others => '0');
   signal ADDR_IN       			: std_logic_vector(7 downto 0) := (others => '0');
   signal NMEA_EN_OUT    			: STD_LOGIC;
   signal NMEA_DATA_OUT  			: STD_LOGIC_VECTOR(7 downto 0);
   signal NMEA_EN_ACK_IN 			: STD_LOGIC;
   signal NEW_TIMESTAMP_EN_OUT   : STD_LOGIC;
	signal TIMESTAMP_DATA_OUT     : STD_LOGIC_VECTOR(31 downto 0);

 	--Outputs
   signal DATA_OUT : std_logic_vector(7 downto 0);

   -- Clock period definitions
   constant CLK_IN_period : time := 10 ns;

   signal TX_OUT        : std_logic := '0';
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: nmea_parser
	PORT MAP (
          CLK_IN          			=> CLK_IN,
          RST_IN          			=> RST_IN,
          NMEA_EN_IN      			=> NMEA_EN_IN,
          NMEA_DATA_IN   			=> NMEA_DATA_IN,
          NMEA_EN_OUT     			=> NMEA_EN_OUT,
          NMEA_DATA_OUT   			=> NMEA_DATA_OUT,
          NMEA_EN_ACK_IN  			=> NMEA_EN_ACK_IN,
			 NEW_TIMESTAMP_EN_OUT   => NEW_TIMESTAMP_EN_OUT,
			 TIMESTAMP_DATA_OUT 		=> TIMESTAMP_DATA_OUT,
          ADDR_IN         			=> ADDR_IN,
          DATA_OUT        			=> DATA_OUT
        );

   uut2: uart
    generic map (
        baud                => 9600,
        clock_frequency     => 100000000
    )
    port map (  
        clock               => CLK_IN,
        reset               => '0',
        data_stream_in      => NMEA_DATA_OUT,
        data_stream_in_stb  => NMEA_EN_OUT,
        data_stream_in_ack  => NMEA_EN_ACK_IN,
        data_stream_out     => open,
        data_stream_out_stb => open,
        tx                  => TX_OUT,
        rx                  => '0'
    );

   -- Clock process definitions
   CLK_IN_process :process
   begin
		CLK_IN <= '0';
		wait for CLK_IN_period/2;
		CLK_IN <= '1';
		wait for CLK_IN_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for CLK_IN_period * 1000;	

--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"56";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4b";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"52";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"43";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"56";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4b";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"52";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"43";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"56";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4b";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"46";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"52";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"43";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"56";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4b";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"56";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"56";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"56";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"52";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"43";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"56";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4b";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"44";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"52";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"43";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"56";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4b";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"43";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"52";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"43";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"53";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"35";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"38";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"45";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"32";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"31";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"36";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"37";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"24";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"50";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"56";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"47";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"33";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"34";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"39";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"54";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4d";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2e";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"4b";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2c";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"2a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"30";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"41";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;
--      NMEA_EN_IN <= '1';
--      NMEA_DATA_IN <= X"0a";
--      wait for CLK_IN_period;
--      NMEA_EN_IN <= '0';
--      wait for CLK_IN_period * 20;

		wait for CLK_IN_period * 10000;
		
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4b";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"43";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"42";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"52";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"43";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4b";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"43";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"52";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"43";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4b";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"43";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"42";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"52";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"43";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4b";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"42";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"52";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"43";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4b";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"52";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"43";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"39";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4b";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"44";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"33";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"52";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"43";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"53";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"38";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"45";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"32";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"36";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"37";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"24";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"50";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"56";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"47";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"31";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"34";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"35";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"54";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4d";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2e";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"4b";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2c";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"41";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"2a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"30";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"44";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;
		NMEA_EN_IN <= '1';
		NMEA_DATA_IN <= X"0a";
		wait for CLK_IN_period;
		NMEA_EN_IN <= '0';
		wait for CLK_IN_period * 20;

    wait for CLK_IN_period * 1000;

    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"24";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"47";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"50";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"5a";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"44";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"41";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"2c";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"30";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"35";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"34";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"32";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"30";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"31";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"2e";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"30";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"30";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"30";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"2c";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"31";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"31";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"2c";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"30";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"32";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"2c";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"32";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"30";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"31";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"36";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"2c";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"2c";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"2a";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"35";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;
    NMEA_EN_IN <= '1';
    NMEA_DATA_IN <= X"33";
    wait for CLK_IN_period;
    NMEA_EN_IN <= '0';
    wait for CLK_IN_period * 20;

      wait;
   end process;

END;
